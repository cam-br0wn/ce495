`ifndef __GLOBALS__
`define __GLOBALS__

// UVM Globals
localparam string THETA_IN_NAME = "../rad.txt";
localparam string COS_OUT_NAME = "../cos_out_uvm.txt";
localparam string SIN_OUT_NAME = "../sin_out_uvm.txt";
localparam string COS_CMP_NAME = "../cos.txt";
localparam string SIN_CMP_NAME = "../sin.txt";
localparam int CLOCK_PERIOD = 10;

`endif
